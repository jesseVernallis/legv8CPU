// bus sizes, in bits
`define COUNTERSIZE     3       // size of the stage counter 
`define BYTESIZE        8       // size of a byte 
`define REGADDRSIZE     5       // size of register address 
`define OPCODESIZE      11      // size of largest opcode 
`define REGDATASIZE     64      // size of a regester in the regester file 
`define INSTRSIZE        32      // size of a instruction 
`define WORDSIZE        32      //size of a word in bits
`define SHAMTSIZE       6       // size of shift amount 
`define SHORTSIZE       26      // size of the largest possible immediate 
