//number of masks used in the control unit
//size of control bus
`define CONTROLSIZE             9

//ID Control Bits
`define REG1ZERO                8
`define REG2LOC                 7
//EX control bits
`define ALUSRC                  6
//DM control bits
`define SETFLAGS                5
`define MEMREAD                 4
`define MEMWRITE                3
//WB control bits               
`define PCTOREG                 2
`define MEMTOREG                1
`define REGWRITE                0

