`include "headers/bus.svh"
`include "headers/sign_extend.svh"

module SignExtend(
input logic[`INSTSIZE-1:0] inst,
input logic[4:0] imm_op,
output logic[`REGDATASIZE-1:0] immediate
);
 
 always_comb begin
	 casex(imm_op)
		//immediate for b type, lsl(2) to word_adress -> byte_adress 
		`IMMOP_B     : immediate = {{36{inst[25]}}, inst[25:0], 2'b0};
		//immediate for cb, lsl(2) to word_adress -> byte_adress 
		`IMMOP_CB    : immediate = {{43{inst[23]}}, inst[23:5], 2'b0};
		`IMMOP_I     : immediate = {52'b0, inst[21:10]};
		`IMMOP_SHIFT : immediate = {58'b0, inst[15:10]};
		`IMMOP_D     : immediate = {{55{inst[20]}}, inst[20:12]};
		 default  : immediate = 64'bx;
	 endcase
 end
endmodule : SignExtend