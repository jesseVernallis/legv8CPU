`define BASE_PATH             "C:/Users/jesse/Desktop/CPU/"
`define INSTUCTION_FILE       {`BASE_PATH, "inst_ram/instructions.txt"}
`define MEM_FILE              {`BASE_PATH, "inst_ram/ram.txt"}