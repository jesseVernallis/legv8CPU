`define IMMCTRL_B        4
`define IMMCTRL_CB       3
`define IMMCTRL_I        2
`define IMMCTRL_SHIFT    1
`define IMMCTRL_D        0

`define IMMOP_B          5'b1xxxx
`define IMMOP_CB         5'b01xxx
`define IMMOP_I          5'b001xx
`define IMMOP_SHIFT      5'b0001x
`define IMMOP_D          5'b00001
`define IMMOP_NONE       5'b00000