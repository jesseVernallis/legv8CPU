
`define MEMPROGSIZE     128     // size of the program memory 
`define MEMDATASIZE     128     // size of the data memory 
`define RAM_FILE                ram file